-- procedure params have direction
-- C <= A+B (matrix)
procedure ADDMATRIX(signal a : in std_logic_vector;
		    signal b : in std_logic_vector;
		    signal c : out std_logic_vector) is
-- local var declarations
begin
	-- sequential statements
end ADDMATRIX;
